`default_nettype none
`timescale 1ns/1ps
/*
this testbench just instantiates the module and makes some convenient wires
that can be driven / tested by the cocotb test.py
*/

// testbench is controlled by test.py
module tb_ticktocktokens ();
    logic [7:0] ui_in;
    logic [7:0] uo_out;
    logic [7:0] uio_in;
    logic [7:0] uio_out;
    logic [7:0] uio_oe;
    logic ena;
    logic clk;
    logic rst_n;

    // this part dumps the trace to a vcd file that can be viewed with GTKWave
    initial begin
        //$dumpfile ("tb.vcd");
        $dumpvars (0, tb_ticktocktokens);
        #1;
    end


    tt_um_jleugeri_ticktocktokens ttt (
        .ui_in(ui_in),
        .uo_out(uo_out),
        .uio_in(uio_in),
        .uio_out(uio_out),
        .uio_oe(uio_oe),
        .ena(ena),
        .clk(clk),
        .rst_n(rst_n)
    );

endmodule : tb_ticktocktokens
